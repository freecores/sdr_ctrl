/*********************************************************************
                                                              
  SDRAM Controller buswidth converter                                  
                                                              
  This file is part of the sdram controller project           
  http://www.opencores.org/cores/sdr_ctrl/                    
                                                              
  Description: SDRAM Controller Buswidth converter

  This module does write/read data transalation between
     application data to SDRAM bus width
                                                              
  To Do:                                                      
    nothing                                                   
                                                              
  Author(s):                                                  
      - Dinesh Annayya, dinesha@opencores.org                 
  Version  :  0.0  - 8th Jan 2012 - Initial structure
              0.2 - 2nd Feb 2012
	         Improved the command pipe structure to accept up-to 4 command of different bank.
                                                              

                                                             
 Copyright (C) 2000 Authors and OPENCORES.ORG                
                                                             
 This source file may be used and distributed without         
 restriction provided that this copyright statement is not    
 removed from the file and that any derivative work contains  
 the original copyright notice and the associated disclaimer. 
                                                              
 This source file is free software; you can redistribute it   
 and/or modify it under the terms of the GNU Lesser General   
 Public License as published by the Free Software Foundation; 
 either version 2.1 of the License, or (at your option) any   
later version.                                               
                                                              
 This source is distributed in the hope that it will be       
 useful, but WITHOUT ANY WARRANTY; without even the implied   
 warranty of MERCHANTABILITY or FITNESS FOR A PARTICULAR      
 PURPOSE.  See the GNU Lesser General Public License for more 
 details.                                                     
                                                              
 You should have received a copy of the GNU Lesser General    
 Public License along with this source; if not, download it   
 from http://www.opencores.org/lgpl.shtml                     
                                                              
*******************************************************************/

`include "sdrc_define.v"
module sdrc_bs_convert (
                    clk,
                    reset_n,
                    sdr_width,

        /* Control Signal from xfr ctrl */
                    x2a_rdstart,
                    x2a_wrstart,
                    x2a_rdlast,
                    x2a_wrlast,
                    app_rd_data_int,
                    app_rd_valid_int,
                    app_wr_data_int,
                    app_wr_en_n_int,
                    app_wr_next_int,

       /* Control Signal from request ctrl */
                    app_req_addr_int,
                    app_req_len_int,
                    app_req_ack_int,
                    app_sdr_req_int,

   /* Control Signal from Bank Ctrl  */
                    app_req_dma_last_int,

   /*  Control Signal from/to to application i/f  */
                    app_req_addr,
                    app_req_len,
                    app_sdr_req,
                    app_req_dma_last,
                    app_req_wr_n,
                    app_req_ack,
                    app_wr_data,
                    app_wr_en_n,
                    app_wr_next,
                    app_rd_data,
                    app_rd_valid
		);
parameter  APP_AW   = 30;  // Application Address Width
parameter  APP_DW   = 32;  // Application Data Width 
parameter  APP_BW   = 4;   // Application Byte Width
parameter  APP_RW   = 9;   // Application Request Width

parameter  SDR_DW   = 16;  // SDR Data Width 
parameter  SDR_BW   = 2;   // SDR Byte Width
   
input                    clk;
input                    reset_n ;
input [1:0]             sdr_width           ; // 2'b00 - 32 Bit SDR, 2'b01 - 16 Bit SDR, 2'b1x - 8 Bit

/* Control Signal from xfr ctrl */
input                    x2a_rdstart; // read start indication
input                    x2a_wrstart; // writ start indication
input                    x2a_rdlast; //  read last burst access
input                    x2a_wrlast; // write last transfer
input [SDR_DW-1:0]       app_rd_data_int;
input                    app_rd_valid_int;
output [SDR_DW-1:0]      app_wr_data_int;
output [SDR_BW-1:0]      app_wr_en_n_int;
input                    app_wr_next_int;

/* Control Signal from request ctrl */
output [APP_AW:0]        app_req_addr_int;
output [APP_RW-1:0]      app_req_len_int; 
input                    app_req_ack_int;
output                   app_sdr_req_int;

/* Control Signal from Bank Ctrl  */
output                   app_req_dma_last_int;


/*  Control Signal from/to to application i/f  */
input [APP_AW-1:0]       app_req_addr;
input  [APP_RW-1:0]      app_req_len ;
input                    app_req_wr_n;
input                    app_sdr_req;
input                    app_req_dma_last;
output                   app_req_dma_last_int;
output                   app_req_ack;

input  [APP_DW-1:0]      app_wr_data;
input  [APP_BW-1:0]      app_wr_en_n;
output                   app_wr_next;

output [APP_DW-1:0]      app_rd_data;
output                   app_rd_valid;

reg [APP_AW:0]           app_req_addr_int;
reg [APP_RW-1:0]         app_req_len_int;

reg                      app_req_dma_last_int;
reg                      app_sdr_req_int;
reg                      app_req_ack;

reg [APP_DW-1:0]         app_rd_data;
reg                      app_rd_valid;
reg [SDR_DW-1:0]         app_wr_data_int;
reg [SDR_BW-1:0]         app_wr_en_n_int;
reg                      app_wr_next;

reg [23:0]               saved_rd_data;
reg [1:0]                rd_xfr_count;
reg [1:0]                wr_xfr_count;


wire                  ok_to_req;                   

assign ok_to_req = ((wr_xfr_count == 0) && (rd_xfr_count == 0));

always @(*) begin
        if(sdr_width == 2'b00) // 32 Bit SDR Mode
          begin
            app_req_addr_int = {1'b0,app_req_addr};
            app_req_len_int = app_req_len;
            app_wr_data_int = app_wr_data;
            app_wr_en_n_int = app_wr_en_n;
            app_req_dma_last_int = app_req_dma_last;
            app_sdr_req_int = app_sdr_req;
            app_wr_next = app_wr_next_int;
            app_rd_data = app_rd_data_int;
            app_rd_valid = app_rd_valid_int;
            app_req_ack = app_req_ack_int;
          end
        else if(sdr_width == 2'b01) // 16 Bit SDR Mode
        begin
           // Changed the address and length to match the 16 bit SDR Mode
            app_req_addr_int = {app_req_addr,1'b0};
            app_req_len_int = {app_req_len,1'b0};
            app_req_dma_last_int = app_req_dma_last;
            //app_sdr_req_int = app_sdr_req && ok_to_req;
            app_sdr_req_int = app_sdr_req ;
            app_req_ack = app_req_ack_int;
            app_wr_next = (app_wr_next_int & wr_xfr_count[0]);
            app_rd_valid = (rd_xfr_count & rd_xfr_count[0]);
            if(wr_xfr_count[0] == 1'b1)
              begin
                app_wr_en_n_int = app_wr_en_n[3:2];
                app_wr_data_int = app_wr_data[31:16];
              end
            else
              begin
                app_wr_en_n_int = app_wr_en_n[1:0];
                app_wr_data_int = app_wr_data[15:0];
              end
            
            app_rd_data = {app_rd_data_int,saved_rd_data[15:0]};
        end else  // 8 Bit SDR Mode
        begin
           // Changed the address and length to match the 16 bit SDR Mode
            app_req_addr_int = {app_req_addr,2'b0};
            app_req_len_int = {app_req_len,2'b0};
            app_req_dma_last_int = app_req_dma_last;
            app_sdr_req_int = app_sdr_req && ok_to_req;
            app_req_ack = app_req_ack_int;
            app_wr_next = (app_wr_next_int & (wr_xfr_count[1:0]== 2'b11));
            app_rd_valid = (rd_xfr_count &   (rd_xfr_count[1:0]== 2'b11));
            if(wr_xfr_count[1:0] == 2'b11)
            begin
                app_wr_en_n_int = app_wr_en_n[3];
                app_wr_data_int = app_wr_data[31:24];
            end
            else if(wr_xfr_count[1:0] == 2'b10)
            begin
                app_wr_en_n_int = app_wr_en_n[2];
                app_wr_data_int = app_wr_data[23:16];
            end
            else if(wr_xfr_count[1:0] == 2'b01)
            begin
                app_wr_en_n_int = app_wr_en_n[1];
                app_wr_data_int = app_wr_data[15:8];
            end
            else begin
                app_wr_en_n_int = app_wr_en_n[0];
                app_wr_data_int = app_wr_data[7:0];
            end
            
            app_rd_data = {app_rd_data_int,saved_rd_data[23:0]};
          end
     end



always @(posedge clk)
  begin
    if(!reset_n)
      begin
        rd_xfr_count    <= 8'b0;
        wr_xfr_count    <= 8'b0;
	saved_rd_data   <= 24'h0;
      end
    else begin

	// During Write Phase
        if(x2a_wrlast) begin
           wr_xfr_count    <= 0;
        end
        else if(app_wr_next_int) begin
           wr_xfr_count <= wr_xfr_count + 1'b1;
        end

	// During Read Phase
        if(x2a_rdlast) begin
           rd_xfr_count    <= 0;
        end
        else if(app_rd_valid_int) begin
           rd_xfr_count   <= rd_xfr_count + 1'b1;
	end

	// Save Previous Data
        if(app_rd_valid_int) begin
	   if(sdr_width == 2'b01) // 16 Bit SDR Mode
	      saved_rd_data[15:0]  <= app_rd_data_int;
            else begin// 8 bit SDR Mode - 
	       if(rd_xfr_count[1:0] == 2'b00)      saved_rd_data[7:0]   <= app_rd_data_int[7:0];
	       else if(rd_xfr_count[1:0] == 2'b01) saved_rd_data[15:8]  <= app_rd_data_int[7:0];
	       else if(rd_xfr_count[1:0] == 2'b10) saved_rd_data[23:16] <= app_rd_data_int[7:0];
	    end
        end
    end
end

endmodule // sdr_bs_convert
